/*
	Anthony De Caria - February 10, 2017
	
	A test Data-stream2
*/

module DS2(index, data);

	/*
		I/O
	*/
	input [5:0] index;
	output reg [109:0] data; 
	
	/*
		Data
	*/
	always @(*)
	begin
		case(index)
			6'b000000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd3000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;		
			end
			6'b000001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd3500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd4000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd4500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd5000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd5500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd6000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd6500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b001000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd7000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd7500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd8000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd8500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd9000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd9500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd10000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd10500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd11000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd11500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd12000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd12500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd13000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b0010101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd13500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b0010110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd14000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd14500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd15000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd15500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd16000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd16500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd17000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd17500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd18000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd18500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd19000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd20000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd20500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd21000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd21500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd22000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd22500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd23000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd23500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd21500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd21500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd21500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd25500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd26000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd26500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd27000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd27500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd28000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd28500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd29000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd29500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd30000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd30500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd31000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd31500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd32000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd32500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd33000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			//change all data below
			6'b111100:
			begin
                data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd215;
                data[23:16] = 8'd215;
                data[31:24] = 8'd100;
                data[47:32] = 16'd33500;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			6'b111101:
			begin
				data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd215;
                data[23:16] = 8'd215;
                data[31:24] = 8'd100;
                data[47:32] = 16'd34000;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			6'b111110:
			begin
				data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd215;
                data[23:16] = 8'd215;
                data[31:24] = 8'd100;
                data[47:32] = 16'd34500;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			6'b111111:
			begin
				data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd215;
                data[23:16] = 8'd215;
                data[31:24] = 8'd100;
                data[47:32] = 16'd35000;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			default:
				data = 110'd0;
		endcase
	end
endmodule

