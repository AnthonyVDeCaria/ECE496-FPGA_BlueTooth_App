/*
	Anthony De Caria - February 9, 2017
	
	A test Data-stream3
*/

module DS3(index, data);

	/*
		I/O
	*/
	input [5:0] index;
	output reg [109:0] data; 
	
	/*
		Data
	*/
	always @(*)
	begin
		case(index)
			6'b000000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd255;
				data[23:16] = 8'd175;
				data[31:24] = 8'd100;
				data[47:32] = 16'd3000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;		
			end
			6'b000001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd254;
				data[23:16] = 8'd176;
				data[31:24] = 8'd100;
				data[47:32] = 16'd3500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd253;
				data[23:16] = 8'd177;
				data[31:24] = 8'd100;
				data[47:32] = 16'd4000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd252;
				data[23:16] = 8'd178;
				data[31:24] = 8'd100;
				data[47:32] = 16'd4500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd251;
				data[23:16] = 8'd179;
				data[31:24] = 8'd100;
				data[47:32] = 16'd5000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd250;
				data[23:16] = 8'd180;
				data[31:24] = 8'd100;
				data[47:32] = 16'd5500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd249;
				data[23:16] = 8'd181;
				data[31:24] = 8'd100;
				data[47:32] = 16'd6000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b000111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd248;
				data[23:16] = 8'd182;
				data[31:24] = 8'd100;
				data[47:32] = 16'd6500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end 
			6'b001000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd247;
				data[23:16] = 8'd183;
				data[31:24] = 8'd100;
				data[47:32] = 16'd7000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd246;
				data[23:16] = 8'd184;
				data[31:24] = 8'd100;
				data[47:32] = 16'd7500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd245;
				data[23:16] = 8'd185;
				data[31:24] = 8'd100;
				data[47:32] = 16'd8000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd244;
				data[23:16] = 8'd186;
				data[31:24] = 8'd100;
				data[47:32] = 16'd8500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd243;
				data[23:16] = 8'd187;
				data[31:24] = 8'd100;
				data[47:32] = 16'd9000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd242;
				data[23:16] = 8'd188;
				data[31:24] = 8'd100;
				data[47:32] = 16'd9500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd241;
				data[23:16] = 8'd189;
				data[31:24] = 8'd100;
				data[47:32] = 16'd10000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b001111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd240;
				data[23:16] = 8'd190;
				data[31:24] = 8'd100;
				data[47:32] = 16'd10500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd239;
				data[23:16] = 8'd191;
				data[31:24] = 8'd100;
				data[47:32] = 16'd11000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd238;
				data[23:16] = 8'd192;
				data[31:24] = 8'd100;
				data[47:32] = 16'd11500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd237;
				data[23:16] = 8'd193;
				data[31:24] = 8'd100;
				data[47:32] = 16'd12000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd236;
				data[23:16] = 8'd194;
				data[31:24] = 8'd100;
				data[47:32] = 16'd12500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd235;
				data[23:16] = 8'd195;
				data[31:24] = 8'd100;
				data[47:32] = 16'd13000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b0010101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd234;
				data[23:16] = 8'd196;
				data[31:24] = 8'd100;
				data[47:32] = 16'd13500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b0010110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd233;
				data[23:16] = 8'd197;
				data[31:24] = 8'd100;
				data[47:32] = 16'd14000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b010111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd232;
				data[23:16] = 8'd198;
				data[31:24] = 8'd100;
				data[47:32] = 16'd14500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd231;
				data[23:16] = 8'd199;
				data[31:24] = 8'd100;
				data[47:32] = 16'd15000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd230;
				data[23:16] = 8'd200;
				data[31:24] = 8'd100;
				data[47:32] = 16'd15500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd229;
				data[23:16] = 8'd201;
				data[31:24] = 8'd100;
				data[47:32] = 16'd16000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd228;
				data[23:16] = 8'd202;
				data[31:24] = 8'd100;
				data[47:32] = 16'd16500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd227;
				data[23:16] = 8'd203;
				data[31:24] = 8'd100;
				data[47:32] = 16'd17000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd226;
				data[23:16] = 8'd204;
				data[31:24] = 8'd100;
				data[47:32] = 16'd17500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd225;
				data[23:16] = 8'd205;
				data[31:24] = 8'd100;
				data[47:32] = 16'd18000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b011111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd224;
				data[23:16] = 8'd206;
				data[31:24] = 8'd100;
				data[47:32] = 16'd18500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd223;
				data[23:16] = 8'd207;
				data[31:24] = 8'd100;
				data[47:32] = 16'd19000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd222;
				data[23:16] = 8'd208;
				data[31:24] = 8'd100;
				data[47:32] = 16'd20000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd221;
				data[23:16] = 8'd209;
				data[31:24] = 8'd100;
				data[47:32] = 16'd20500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd220;
				data[23:16] = 8'd210;
				data[31:24] = 8'd100;
				data[47:32] = 16'd21000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd219;
				data[23:16] = 8'd211;
				data[31:24] = 8'd100;
				data[47:32] = 16'd21500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd218;
				data[23:16] = 8'd212;
				data[31:24] = 8'd100;
				data[47:32] = 16'd22000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd217;
				data[23:16] = 8'd213;
				data[31:24] = 8'd100;
				data[47:32] = 16'd22500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b100111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd216;
				data[23:16] = 8'd214;
				data[31:24] = 8'd100;
				data[47:32] = 16'd23000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd215;
				data[23:16] = 8'd215;
				data[31:24] = 8'd100;
				data[47:32] = 16'd23500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd214;
				data[23:16] = 8'd216;
				data[31:24] = 8'd100;
				data[47:32] = 16'd24000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd213;
				data[23:16] = 8'd217;
				data[31:24] = 8'd100;
				data[47:32] = 16'd24500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd212;
				data[23:16] = 8'd218;
				data[31:24] = 8'd100;
				data[47:32] = 16'd25000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd211;
				data[23:16] = 8'd219;
				data[31:24] = 8'd100;
				data[47:32] = 16'd25500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd210;
				data[23:16] = 8'd220;
				data[31:24] = 8'd100;
				data[47:32] = 16'd26000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd209;
				data[23:16] = 8'd221;
				data[31:24] = 8'd100;
				data[47:32] = 16'd26500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b101111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd208;
				data[23:16] = 8'd222;
				data[31:24] = 8'd100;
				data[47:32] = 16'd27000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd207;
				data[23:16] = 8'd223;
				data[31:24] = 8'd100;
				data[47:32] = 16'd27500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd206;
				data[23:16] = 8'd224;
				data[31:24] = 8'd100;
				data[47:32] = 16'd28000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd205;
				data[23:16] = 8'd225;
				data[31:24] = 8'd100;
				data[47:32] = 16'd28500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd204;
				data[23:16] = 8'd226;
				data[31:24] = 8'd100;
				data[47:32] = 16'd29000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110100:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd203;
				data[23:16] = 8'd227;
				data[31:24] = 8'd100;
				data[47:32] = 16'd29500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110101:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd202;
				data[23:16] = 8'd228;
				data[31:24] = 8'd100;
				data[47:32] = 16'd30000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110110:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd201;
				data[23:16] = 8'd229;
				data[31:24] = 8'd100;
				data[47:32] = 16'd30500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b110111:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd200;
				data[23:16] = 8'd230;
				data[31:24] = 8'd100;
				data[47:32] = 16'd31000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111000:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd199;
				data[23:16] = 8'd231;
				data[31:24] = 8'd100;
				data[47:32] = 16'd31500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111001:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd198;
				data[23:16] = 8'd232;
				data[31:24] = 8'd100;
				data[47:32] = 16'd32000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111010:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd1;
				data[15:8] = 8'd197;
				data[23:16] = 8'd233;
				data[31:24] = 8'd100;
				data[47:32] = 16'd32500;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			6'b111011:
			begin
				data[6:0] = 7'd77;
				data[7] = 1'd0;
				data[15:8] = 8'd196;
				data[23:16] = 8'd234;
				data[31:24] = 8'd100;
				data[47:32] = 16'd33000;
				data[55:48] = 8'd239;
				data[63:56] = 8'd17;
				data[79:64] = 16'd0;
				data[85:80] = 6'd1;
				data[109:86] = 24'd4272433;
			end
			//change all data below
			6'b111100:
			begin
                data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd195;
                data[23:16] = 8'd235;
                data[31:24] = 8'd100;
                data[47:32] = 16'd33500;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			6'b111101:
			begin
				data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd194;
                data[23:16] = 8'd236;
                data[31:24] = 8'd100;
                data[47:32] = 16'd34000;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			6'b111110:
			begin
				data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd193;
                data[23:16] = 8'd237;
                data[31:24] = 8'd100;
                data[47:32] = 16'd34500;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			6'b111111:
			begin
				data[6:0] = 7'd77;
                data[7] = 1'd0;
                data[15:8] = 8'd192;
                data[23:16] = 8'd238;
                data[31:24] = 8'd100;
                data[47:32] = 16'd35000;
                data[55:48] = 8'd239;
                data[63:56] = 8'd17;
                data[79:64] = 16'd0;
                data[85:80] = 6'd1;
                data[109:86] = 24'd4272433;
			end
			default:
				data = 110'd0;
		endcase
	end
endmodule

